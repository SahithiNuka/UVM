package d_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "d_trans.sv"
	`include "d_cfg.sv"
	`include "d_driver.sv"
	`include "d_monitor.sv"
	`include "d_seqr.sv"
	`include "d_agent.sv"
	`include "d_seqs.sv"
	`include "d_sb.sv"
	`include "d_env.sv"
	`include "d_test.sv"

endpackage
