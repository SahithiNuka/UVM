package p_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "p_trans.sv"
	`include "p_cfg.sv"
	`include "p_driver.sv"
	`include "p_monitor.sv"
	`include "p_seqr.sv"
	`include "p_agent.sv"
	`include "p_seq.sv"
	`include "p_sb.sv"
	`include "p_env.sv"
	`include "p_test.sv"

endpackage
