interface inf();
	logic [7:0]in;
	logic [2:0]out;
	
	modport MP(input out, output in);
endinterface